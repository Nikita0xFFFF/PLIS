package crc_pkg;
  localparam  write_crc8 = 32'd0;
  localparam  read_crc8 = 32'd4;
  localparam  write_crc15 = 32'd8;
  localparam  read_crc15 = 32'd12;
  
endpackage : crc_pkg
